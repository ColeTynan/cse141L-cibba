// Module Name:    InstFetch 
// Project Name:   CSE141L
//
// Revision Fall 2020
// Based on SystemVerilog source code provided by John Eldon
// Comment:
// This module does not actually fetch the actual code
// It is responsible for providing which line number will be read next


	 
module InstFetch(Reset,Start,clk,branch_abs,branch_rel_en,ALU_flag,target,prog_ctr);

  input              Reset,			   // reset, init, etc. -- force PC to 0 
                     Start,			   // begin next program in series
                     clk,			      // PC can change on pos. edges only
                     branch_abs,	       // jump unconditionally to target value	   
                     branch_rel_en,	   // jump conditionally to target + PC
                     ALU_flag;		   // flag from ALU, e.g. Zero, Carry, Overflow, Negative (from ARM)
  input       [9:0] target;		      // jump ... "how high?"
  output reg[9:0] prog_ctr ;            // the program counter register itself
  
  
  //// program counter can clear to 0, increment, or jump
	always
	begin 
		if(Reset)
		  prog_ctr <= 0;				        // for first program; want different value for 2nd or 3rd
		else if(Start)						     // hold while start asserted; commence when released
		  prog_ctr <= prog_ctr;
		else if(branch_abs)	              // unconditional absolute jump
		  prog_ctr <= target;
		else if(branch_rel_en && ALU_flag)   // conditional relative jump
		  prog_ctr <= target + prog_ctr;
		else
		  prog_ctr <= prog_ctr+'b1; 	        // default increment (no need for ARM/MIPS +4. Pop quiz: why?)
	end


endmodule

/* Note about Start: if your programs are spread out, with a gap in your machine code listing, you will want 
to make Start cause an appropriate jump. If your programs are packed sequentially, such that program 2 begins 
right after Program 1 ends, then you won't need to do anything special here. 
*/